
module and_power (input i1, i2, i3, i4, clk,
                  output out);

    assign out = i1 & i2 & i3 & i4;

endmodule


