
module simple (input  [1:0] x, 
               output [1:0] y);
    assign y = ~x;
endmodule




